module pin

#define pin__write(PIN_NAME, VALUE)   digitawrite(PIN_NAME, VALUE)