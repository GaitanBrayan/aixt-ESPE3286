module pin

<<<<<<< HEAD
#define pin__out OUTPUT

#define pin__in INPUT_PULLUP
=======
#define pin__output		OUTPUT
#define pin__input		INPUT
#define pin__in_pullup	INPUT_PULLUP

fn init() {

}
>>>>>>> 2d8f797db8c3c5c757c2f3c7abe22d9bbd8f42fb
