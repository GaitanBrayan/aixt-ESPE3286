module adc

#define adc__write(PIN_NAME, MODE)   analogWrite(PIN_NAME, MODE)