module time

#define time__sleep_ms(MS)  delay(MS)