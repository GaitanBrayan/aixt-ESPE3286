module pin

#define pin__mode(PIN_NAME, MODE)    pinMode(PIN_NAME, MODE)