<<<<<<< HEAD
module time 
=======
module time


fn init() {

}
>>>>>>> 2d8f797db8c3c5c757c2f3c7abe22d9bbd8f42fb
