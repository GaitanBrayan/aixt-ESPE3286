module time 