module port