module port
define port__read(PORT_NAME)  PORT ## PORT_NAME