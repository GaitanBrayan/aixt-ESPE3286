module port

define port__write(PORT_NAME, VALUE)	LAT ## PORT_NAME = VALUE