module pin

<<<<<<< HEAD
#define pin__setup(PIN_NAME, MODE)   digitalSETUP(PIN_NAME, MODE)
=======
#define pin__setup(PIN_NAME, MODE)    pinMode(PIN_NAME, MODE)
>>>>>>> 2d8f797db8c3c5c757c2f3c7abe22d9bbd8f42fb
