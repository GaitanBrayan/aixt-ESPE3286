module uart

#define uart0__setup_1(BAUD_RATE)   Serial.begin(BAUD_RATE).,