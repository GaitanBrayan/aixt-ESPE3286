module pin

<<<<<<< HEAD
#define pin__write(PIN_NAME, VALUE)   digitawrite(PIN_NAME, VALUE)
=======
#define pin__write(PIN_NAME, VALUE)   digitalWrite(PIN_NAME, VALUE)
>>>>>>> 2d8f797db8c3c5c757c2f3c7abe22d9bbd8f42fb
