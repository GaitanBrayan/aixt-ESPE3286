module port

define port__setup(PORT_NAME, VALUE)   TRIS ## PORT_NAME = VALUE