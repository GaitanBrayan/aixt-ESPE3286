module pin

#define pin__setup(PIN_NAME, MODE)   digitalSETUP(PIN_NAME, MODE)