module time

#define time__sleep_us(US)  delayMicroseconds(US)